library verilog;
use verilog.vl_types.all;
entity RTLDesign_vlg_vec_tst is
end RTLDesign_vlg_vec_tst;
